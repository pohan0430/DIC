
module PATTERN	(
	// output
    IFM_0, IFM_1, IFM_2, IFM_3,
	INW_0, INW_1, INW_2, INW_3,
	//input
	Output,

);

//------------------------------
//	I/O Pors
//------------------------------
output reg [3:0] IFM_0, IFM_1, IFM_2, IFM_3;
output reg [3:0] INW_0, INW_1, INW_2, INW_3;

input wire[9:0]Output;
reg [9:0]Golden_Output;

integer i, j;
parameter PAT_NUM=1000;

reg figure;

initial begin
	IFM_0='d0; IFM_1='d0; IFM_2='d0; IFM_3='d0;
	INW_0='d0; INW_1='d0; INW_2='d0; INW_3='d0;
	Golden_Output = 'd0;	
	
	#100;

	for(i=0;i<PAT_NUM;i=i+1)begin
		IFM_0=$urandom_range(15,0); IFM_1=$urandom_range(15,0); 
		IFM_2=$urandom_range(15,0); IFM_3=$urandom_range(15,0); 
		INW_0=$urandom_range(15,0); INW_1=$urandom_range(15,0); 
		INW_2=$urandom_range(15,0); INW_3=$urandom_range(15,0); 
		Golden_Output=IFM_0*INW_0+IFM_1*INW_1+IFM_2*INW_2+IFM_3*INW_3;
		#100;
		check_ans_task;
	end
	`ifdef RTL
	PASS_RTL;
	`endif	
	`ifdef GATE
	PASS_GATE;
	`endif
end



task check_ans_task; begin
	//#(5)
		if(Output !== Golden_Output) begin
					$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
					$display ("                                                                        OUTPUT FAIL!                                                               ");
					$display ("                                                                   PATTERN NO.%4d                                                           ",j);
					$display ("                                                     Ans(OUT): %d,  Your output : %d  at %8t                                              ",Golden_Output,Output,$time);
					$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
					$finish;
		end	
end endtask





task PASS_RTL;begin
$display("                                                                                        \033[0;40;34m```....``\033[0;40;37m                                                                                   ");
$display("                                                                             \033[0;40;34m`-:/+osyyhhhhhhhhhhhhyso/:.`\033[0;40;37m                                                                           ");
$display("                                                                       \033[0;40;34m.:/oyhhhhyyyyyyyyyyyyyyyyyyyyyyyyhyo/:.\033[0;40;37m                                                                      ");
$display("                                                                  \033[0;40;34m.:+shhyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyhys/-`\033[0;40;37m                                                                 ");
$display("                                                              \033[0;40;34m-/oyhyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyys/-\033[0;40;37m                                                              ");
$display("                                                          \033[0;40;34m./shhyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyo:`\033[0;40;37m                                                          ");
$display("                                                       \033[0;40;34m./shyyyyyyyyyyyyyyyyyyyyyyysso++/::--......-://+osyyyyyyyyyyyyyyyyys:`\033[0;40;37m                                                       ");
$display("                                                    \033[0;40;34m`:syyyyyyyyyyyyyyyyyyyyyso+/-.```                  ``.-:+ossyyyyyyyyyyyyyo:`\033[0;40;37m                                                    ");
$display("                                                  \033[0;40;34m-os+/yyyyyyyyyyyyyyyss+/-.`                                 ``-:+osyyyyyyys/+so-\033[0;40;37m                                                  ");
$display("                                               \033[0;40;34m`:so/:-/syyyyyyyyyyso/:.`                                           ``-/+syyyyo::/os/`\033[0;40;37m                                               ");
$display("                                             \033[0;40;34m`/so:---:syyyyyyyys+:``\033[0;40;37m                `.-::::::::::::::---.`              \033[0;40;34m`-/osys+:::+so-\033[0;40;37m   ");
$display("                                           \033[0;40;34m`/so:---:+syyyyyso/.`\033[0;40;37m             `.-:///:-.`````       ````..-:/::-.`          \033[0;40;34m`.:+ssssosyhs-\033[0;40;37m   ");
$display("                                         \033[0;40;34m`/yy+///+ossyyyyo/.`\033[0;40;37m            .-://-.``      .o+-      `+o/`     ``.-:/:-.          \033[0;40;34m`-+syyyyyhs:\033[0;40;37m    ");
$display("                                        \033[0;40;34m:yhyyysssyyyyys+-`\033[0;40;37m           `-:/:.`   -/.     :o:-++.   :o/.:o:`   -+o:  `.-/:-.         \033[0;40;34m.:osyyyyhs:\033[0;40;37m    ");
$display("                                      \033[0;40;34m.ohyyyyyyyyyyys/.\033[0;40;37m           .://-.     `++:++:..o/.```-+/-o/.```.:o::o/-.++`    `-:/:-        \033[0;40;34m`.+syyyyhs-\033[0;40;37m    ");
$display("                                     \033[0;40;34m/yyyyyyyyyyyys/.\033[0;40;37m          `://.``++/:` .o/.```-:/-```````-/-````````::.````:o- `-+++``-/:-`       \033[0;40;34m./syyyyho.\033[0;40;37m    ");
$display("                                   \033[0;40;34m.shyyyyyyyyyys+.\033[0;40;37m         `-//-`  .o:.-:/+o-`````.`````````````````````````````.+++:../o.  `-//-`      \033[0;40;34m`:oyyyhy/\033[0;40;37m    ");
$display("                                  \033[0;40;34m:yyyyyyyyyyyso-\033[0;40;37m         .:+/+:.  :+.````````````.:.``````````````````````````````.`````-o:  ./:-/:.      \033[0;40;34m`:syyyhs.\033[0;40;37m    ");
$display("                                \033[0;40;34m`+hyyyyyyyyyys:`\033[0;40;37m        -//..o::/++/``````````````-/:```````````````````````````.`````````.+++/-o: .:/-`     \033[0;40;34m`/syyyh:\033[0;40;37m    ");
$display("                               \033[0;40;34m`ohyyyyyyyyys/`\033[0;40;37m       `-+/. :o-````.```````````.```-//-`..```````````````````````+.``````````.````+/` `-//.     \033[0;40;34m.+syyh+`\033[0;40;37m    ");
$display("                              \033[0;40;34m.shyyyyyyyys+.\033[0;40;37m       `-+o:``++``````````````````:.``-///.--```````````````````````:s````````````````/o../:.//.     \033[0;40;34m-oyyhs.\033[0;40;37m    ");
$display("                             \033[0;40;34m.yhyyyyyyyys-\033[0;40;37m        -+:/o:/+:``````````````````/+-``-///:-:```````````````````````.h/````````````````-+/-/o.`//.    \033[0;40;34m`+syhy.\033[0;40;37m    ");
$display("                            \033[0;40;34m.yyyyyyyyys+`\033[0;40;37m       -+/`/o.``````````````````````oo:``-//////-```````````````````````y+-````````.```````````-o/`.+/`    \033[0;40;34m:syhh.\033[0;40;37m    ");
$display("                           \033[0;40;34m.yhyyyyyyys/`\033[0;40;37m      `++``++````````````..``````````ys/-`-//////:```````````````````````h.o`````````-.```````````:o/++o-    \033[0;40;34m.oyhh.\033[0;40;37m    ");
$display("                          \033[0;40;34m`yhyyyyyyys:\033[0;40;37m       :o++/+/```````````./.``````````-oy/:`.///////.``````````````````````h`+-```````/`--.```````````:``.+/`   \033[0;40;34m`oyhy.\033[0;40;37m    ");
$display("                         \033[0;40;34m`shyyyyyyys:\033[0;40;37m      .o+..`..```````````-o-..`````````o.o+/-`///////:````````````-````````.h -o```````o/`./+``````````````.:o`   \033[0;40;34m`oyhy`\033[0;40;37m    ");
$display("                         \033[0;40;34mohyyyyyyys:\033[0;40;37m      :o:.```````````````:o:-.``./.````:+`:h//.:///////-```````````s````````:y-.y```````/-+`./o```````````````-o.   \033[0;40;34m`oyho\033[0;40;37m    ");
$display("                        \033[0;40;34m/hyyyyyyys:\033[0;40;37m     `+o..```````````````-s/-.``:o+````.s::.oo/:-////////``````````-s:```````o:`-y:.`````-/.o`-+o```````````````-o-   \033[0;40;34m.syd/\033[0;40;37m    ");
$display("                       \033[0;40;34m-dyyyyyyyy/\033[0;40;37m     `o/..```````````````.s/:.`:/:+```.:s:`  `s//:////////:`````````o-+```````y`  +/-::-.`.o -o`-+o```````````````.s.   \033[0;40;34m:syh.\033[0;40;37m    ");
$display("                      \033[0;40;34m`yhyyyyyyyo\033[0;40;37m     `s/.`````````````````o+:-:/..o-::::s-     .s///////////-```````-h`o``````//   /:```--:/s.`//`:o+```````````````.s.   \033[0;40;34moyhs\033[0;40;37m    ");
$display("                      \033[0;40;34m+hyyyyyyys.\033[0;40;37m    `s:.`````````````````-y/++:-/o:-.`.+.       ./+++++////++:.----:o/ o--...-+`   //------:+..`s.-/s-```````````````-o`  \033[0;40;34m.syd:\033[0;40;37m    ");
$display("                     \033[0;40;34m.dyyyyyyys:\033[0;40;37m    `s:.``````````````````os/.`` /////:-`          ``..---::::----..``  `......     `..-.--..`   .::+oy````````````````:+   \033[0;40;34m/yhh/`\033[0;40;37m    ");
$display("                     \033[0;40;34msdyyyyyyyo\033[0;40;37m     o/.``````````:````````y`                                                                          +/````````````````+:  \033[0;40;34m`sydhy-\033[0;40;37m    ");
$display("                    \033[0;40;34m:hyyyyyyys.\033[0;40;37m    /o.```````````+-``````.s                                                                           .y```````:````````.y   \033[0;40;34m/yhhyho.\033[0;40;37m    ");
$display("                  \033[0;40;34m.ohyyyyyyyy+\033[0;40;37m    .y.````````````:+``````:o                                                                            y.`````-/`````````y-  \033[0;40;34m.sydyyyh/\033[0;40;37m    ");
$display("                 \033[0;40;34m/hyyyyyyyyyy-\033[0;40;37m    o/.`````````````y.`````:+                                                                            +:`````o.`````````o+   \033[0;40;34moydyyyyhs.\033[0;40;37m    ");
$display("              \033[0;40;34m`shyyyyyyyyyyo\033[0;40;37m    .y.``````````````:s`````:o`ooooooooo+++//::-.`````                              ```.--:::///++++++/-  //````.s``````````/s   \033[0;40;34m/yhhyyyyyh:\033[0;40;37m   ");
$display("              \033[0;40;34m-hhyyyyyyyyyyy/\033[0;40;37m    +o-```````````````++````-s-ddddddddddddddddddddhyy/                            /yhdddddddddddhhhhhho  /+````s-``````````-y   \033[0;40;34m.yydyyyyyyh+\033[0;40;37m    ");
$display("             \033[0;40;34m:hyyyyyyyyyyyyy-\033[0;40;37m    y//````````````````++```.y ```````....--::/+hdddddo                            /hdddh+-.`````         //```o:```````````.h`  \033[0;40;34m`sydyyyyyyyho`\033[0;40;37m    ");
$display("            \033[0;40;34m/dyyyyyyyyyyyyys`\033[0;40;37m   .s:+`````````````````/o.``s`             `/sdddds/`               `      `        -/sdddho:`           o-``o:`````````````h`   \033[0;40;34moyhhyyyyyyyhs\033[0;40;37m    ");
$display("           \033[0;40;34m/dyyyyyyyyyyyyyyo\033[0;40;37m    :+/+``````````````````.o:`//          `/sdddho:`           `    ``      `      `     `-+ydddy/.       `y`-o-`````````-````y.   \033[0;40;34m/yhhyyyyyyyyho\033[0;40;37m    ");
$display("          \033[0;40;34m/dyyyyyyyyyyyyyyy+\033[0;40;37m    //+/````````````````````++-o       `:sdddho:`                  ``      `      `          ./sdddy/.    -+/o``````````::````o/   \033[0;40;34m:yhhyyyyyyyyyh+\033[0;40;37m    ");
$display("         \033[0;40;34m:dyyyyyyyyyyyyyyyy/\033[0;40;37m    +/s-````````````````````:/`-`   `-ohddds:`               .-:-.`      ``  `-::::.            `:ohddy/` :-`o``````````s`````-y   \033[0;40;34m:yhdyyyyyyyyyyd-\033[0;40;37m    ");
$display("        \033[0;40;34m-dyyyyyyyyyyyyyyyyy/\033[0;40;37m    /oy``````````````````````y`   -+hddds/`               `////.-+//+:`    -+s:./:.oo`             `-ohdo   `s`````````/+``````y:  \033[0;40;34m:yydyyyyyyyyyyyy`\033[0;40;37m    ");
$display("       \033[0;40;34m`yhyyyyyyyyyyyyyyyyy+\033[0;40;37m    -d+``````````````````````+:  -hddy/.`                 o++/://:/+:/o/:/+++::/::/::s`         \033[0;40;31m```````.`\033[0;40;37m   -o````````-s```````-y` \033[0;40;34m/yhdyyyyyyyyyyyh/\033[0;40;37m    ");
$display("       \033[0;40;34m+dyyyyyyyyyyyyyyyyyyo\033[0;40;37m    `h.``````````````````````.y`  \033[0;40;31m-/.````````````````\033[0;40;37m    -o::::::::::::::::::::::::::y-   \033[0;40;31m``````````````````\033[0;40;37ms-```````-s.````````+s \033[0;40;34moyhhoyhyyyyyyyyh+\033[0;40;37m    ");
$display("      \033[0;40;34m`dyyyyyyyyyyyyyyyyyyys\033[0;40;37m    ++````````````````````````:s` \033[0;40;31m``````````````````````\033[0;40;37m :+::::::::::::::::::::::::::y.  \033[0;40;31m``````````````````\033[0;40;37m:o```````/o```````````oos\033[0;40;34msdo `.:+syhyyhy.\033[0;40;37m    ");
$display("      \033[0;40;34m-dyyyyyyyyyyyyyyhyyyyy.\033[0;40;37m  -s``````````````````````````/o\033[0;40;31m```````````````````````\033[0;40;37m `s::::::::::++/:-:/+/::::::/o   \033[0;40;31m`````````````````\033[0;40;37m-y.`````.o/``./:````````+h\033[0;40;34myd-      ``..``\033[0;40;37m     ");
$display("       \033[0;40;34moyhhhhyyyso+/:-hyyyyy/\033[0;40;37m .y.`````````.-`````--`````````+o\033[0;40;31m`````````````````````\033[0;40;37m   -++/::///+/.`     `://////:`     \033[0;40;31m``````````````\033[0;40;37m-s-`````/+.`````-//:``````:yh`\033[0;40;37m                 ");
$display("        \033[0;40;34m````````      ohyyyys\033[0;40;37m.s-`````````:+```````-/-````````/o.\033[0;40;31m````````````````\033[0;40;37m       ``-:--.``           `````\033[0;40;37m                    -o.```./+-`````````.-s+:-```.+o.\033[0;40;37m                ");
$display("                      \033[0;40;34m.dyyyyy\033[0;40;37ms.````````:+:``````````:+:.``````-o-\033[0;40;31m````````\033[0;40;37m                                                         `//```:+/.`````````````h`.:so/:--//-`\033[0;40;37m             ");
$display("                       \033[0;40;34mshyy\033[0;40;37myo.``````.:s:``````````````-//:.````.+/`                                                             `-/-.-:sh:`.````````````:s  `syd:-://++-\033[0;40;37m            ");
$display("                       -dys:`````.://-o.`````````````.-``-/++:-.`-/:`                                                           `.````/h:`.:````````````s/  \033[0;40;34m+yho\033[0;40;37m                    ");
$display("                       .o/.`.-:+/:.`  -+``````````````:.````+/-:///+o/-`                                                            `oy-``:.```````````.h` \033[0;40;34m-syy`\033[0;40;37m                    ");
$display("                    .//:+sssyyy:      y.`````````````.:````.s`  ```````                                                           -y+.``-:````````````o+ `\033[0;40;34msyh.\033[0;40;37m                     ");
$display("                         \033[0;40;34m`yhyyyys-\033[0;40;37m     :o``````````````--````sh/.                                                                .os:```-/.``.````````:y``\033[0;40;34m+yh-\033[0;40;37m                      ");
$display("                          \033[0;40;34m`shyyyys-\033[0;40;37m     o:``````````.```:.```-hyy+.                                                            .+s/````-/:``-.```````.y- \033[0;40;34m/yy-\033[0;40;37m                       ");
$display("                          \033[0;40;34m `ohyyyys-\033[0;40;37m    `s-`````````--``.:-```+o-oys:.                                                      `-+o:.````-/:``--````````s+`\033[0;40;34m/hs.\033[0;40;37m                        ");
$display("                          \033[0;40;34m   :yyyyys:\033[0;40;37m    .s-`````````:-``-/-```s: `:oso:`      ``                                  `     `-/s/-``````://-`-:`..`````oo.\033[0;40;34m+y/`\033[0;40;37m                         ");
$display("                          \033[0;40;34m    .+yyyys/`\033[0;40;37m   .o:`````````::.`-/-``.s:   .:oso:.``:++:`     .:`      ..       ./.    `/+/..-/+:-s``````.://:.:/.`o.````oo:\033[0;40;34mso.\033[0;40;37m                           ");
$display("                          \033[0;40;34m      ./yyyyo.\033[0;40;37m   `+/````````.::.`-/:.`.s:     `-+ooso-.:+-``-/:-o:   `/+++.   `:o-+/``:o/-+o:-.  /:`.-``.:///-:/-`/y```.sso\033[0;40;34ms-\033[0;40;37m                             ");
$display("                          \033[0;40;34m        `syyys/`\033[0;40;37m   /+.```-/```:/:.-//-..s:        `-/+ooohss/-```++.:+-  -+/.-o/..-+o/+:-.`     .o`:+/`-////://-`/s+``-yhs:\033[0;40;34m`\033[0;40;37m                              ");
$display("                                   o/\033[0;40;34m-+yhs:`\033[0;40;37m  .+/```s+.``-:/:://:-.o+`           `.-:/++++++oss/::::/sso/-...``          `o:/-+::///////:.//o.`+hh-                                 ");
$display("                                   o:`\033[0;40;34m`.:oys:`\033[0;40;37m  -+-`-o+:``.://////:-/o.                     `````  ```./+.              .so/``y////////:-+://-o//o                                  ");
$display("                                   y-```\033[0;40;34m``.:oo+:\033[0;40;37m.`:/-:+:+/.`-://////:/s/`                      `..`     :y            `:s+.  +o//+o///:+s+ss++.`/o                                  ");
$display("                                  `h````````\033[0;40;34m``-/+o\033[0;40;37m+//+/o--/+:.-:///os+/oo:`                  `+///++    .y            .-`   :s/+os+//oyyoyy/.```/o                                  ");
$display("                                  :o``````````````-/+osyho--:/+/:///+soo+oo:`                `++/++/   -s-                 -s+so+o/+/:..--``````-y                                  ");
$display("                                  s:```````````````....-:/+oooossyyysssso:-:.                  ``.``.:+/.           ```.-:+yssos+::``````````````h.                                 ");
$display("                                 -y```````````````............--:://+++oosyo+///::::::::://++++++++oss+///::::::/+oo++++//:-.......``````````````o+                                 ");
$display("                                 s:```````````````.......................:y```..---------..+:.```   .+` ``````````-s................`````````````-h`                                ");
$display("                                /s```````````````........................:hs/.`             :/.````.o`            `y................``````````````o/                                ");
$display("                               .y.````..````````...............:........\033[0;40;34mohyyyyso/-``\033[0;40;37m       `//y++++y:/`      \033[0;40;34m`.:+oyy/\033[0;40;37m....--..........`````````````.h.                               ");
$display("                              `s/````:s`````````.............../......-\033[0;40;34myyyyyyyyyyyyso+:.``\033[0;40;37m  ..-+++o/..  \033[0;40;34m`.:+oyyyyyyyho\033[0;40;37m..../..........``````````-```:y`                              ");
$display("                              o+````+oo````````../............+-.....:\033[0;40;34myyyyyyyyyyyyyyyhooss+::o--s+o`:/:oys+oyyyyyyyyyys-\033[0;40;37m..::..........`````````:+```+o                              ");
$display("                             +o```-o-+/```````../o...........:+.....:\033[0;40;34mhyyyyyyyyyyyyyyyy\033[0;40;37m::\033[0;40;34myyyyyyo::h-:oyyyyy\033[0;40;37m::\033[0;40;34myyyyyyyyyyyy\033[0;40;37m-..o...........-````````os.``o+                             ");
$display("                            +o``.++` y.``````..:h-...........s-....:\033[0;40;34mhyyyyyyyyyyyyyyyh+\033[0;40;37m:\033[0;40;34m+hyyyyyyyyhydhhyyyh+\033[0;40;37m:\033[0;40;34m/hyyyyyyyyyyy\033[0;40;37m-.//..........+-````````yo/``o+                            ");
$display("                          `s/`.+o.  :o``````..-ho...........+/....-\033[0;40;34mhyyyyyyyyyyyyyyyyy\033[0;40;37m::\033[0;40;34myyyyyyhhhhdhhhyyyyyy\033[0;40;37m::\033[0;40;34msyyyyyyyyyyyy\033[0;40;37m..+-..........o-```````-s:o-`++                           ");
$display("                         -s--++.    y-`````..-ys-........../o.....\033[0;40;34myyyyyyyyyyyyyyyyyyo\033[0;40;37m::\033[0;40;34mhyyyyyydhhyyyyyyyyyh/\033[0;40;37m:\033[0;40;34m/hyyyyyyyyyyhs\033[0;40;37m.:/-.........-y:```````/+`/o./s`                         ");
$display("                       .oo++/`     :o`````..-y:o..........:+:....\033[0;40;34m+hyyyyyyyyhyyyyyyyh/\033[0;40;37m:\033[0;40;34m+hyyyyyyyyyyyyyyyyyyho\033[0;40;37m::\033[0;40;34myyyyhyyyyyyyh\033[0;40;37m+.//..........:h/```````+/ `+o/s:                        ");
$display("                     .oh+/.       `y.```...:y.s-.........-/+....-\033[0;40;34mhyyyyyyyyyhyyyyyyyh\033[0;40;37m::\033[0;40;34mohyyyyyyyyyyyyyyyyyyyy\033[0;40;37m::\033[0;40;34moyyyhyyyyyyyyh\033[0;40;37m-.//..........+y+```````o:  `/+so.                      ");
$display("                   `--`           s:```.../s`//.........-/+.....\033[0;40;34msyyyyyyyyyyhyyyyyyyy\033[0;40;37m::\033[0;40;34msyyyyyyyyyyyyyyyyyyyyh/\033[0;40;37m:\033[0;40;34m/hyyyhyyyyyyyyy\033[0;40;37m.:-/..........+oo-``````o/    `:+/`                    ");

$display ("----------------------------------------------------------------------------------------------------------------------");
$display ("                                                  Congratulations!                						            ");
$display ("----------------------------------------------------------------------------------------------------------------------");
$finish;	
end endtask

task PASS_GATE;begin
  $display("                                                             \033[33m                                                                             ");        
  $display("                                                             /NN.                                                                           ");        
  $display("                                                            sMMM+                                                                           ");        
  $display("                                                           sMMMMy                                                                           ");        
  $display(" oNNmhs+:-                                                oMMMMMh                                                                           ");        
  $display("  /mMMMMMNNd/:-                                          :+smMMMh                                                                           ");        
  $display("   .sNMMMMMN::://:-                                     .o--:sNMy                                                                           ");        
  $display("     -yNMMMM:----::/:-.                                 o:----/mo                                                                           ");        
  $display("       -yNMMo--------://:.                             -+------+/                                                                           ");        
  $display("         .omd/::--------://:                           o-------o.                                                                           ");        
  $display("           `/+o+//::-------:+:                        .+-------y                                                                            ");        
  $display("              .:+++//::------:+/.---------.           +:------/+                                                                            ");        
  $display("                 `-/+++/::----:/:::::::::::://:-.     o------:s.          \033[30m:::::----.           -::::.          `-:////:-`     `.:////:-.    \033[33m");        
  $display("                    `.:///+/------------------:::/:- `o-----:/o          \033[31m NNNNNNNNNNds-        NNNNNN        .smNMMMMMMNy   .smNNMMMMMNh    \033[33m");        
  $display("                         :+:----------------------::/:s-----/s.          \033[31m MMMMo++sdMMMN-      mMMmMMMs      -NMMMh+///oys   mMMMdo///oyy    \033[33m");        
  $display("                        :/---------------------------:++:--/++           \033[32m MMMM.    mMMMy     yMMM:dMMM/     +MMMM:         :MMMM+           \033[33m");        
  $display("                       :/---///:-----------------------::-/+o`           \033[32m MMMM.    NMMMo    +MMMs -NMMm.    .mMMMNdo:.     `dMMMNds/-       \033[33m");        
  $display("                      -+--/dNs-o/------------------------:+o`            \033[36m MMMMyyyhNMMNy    -NMMm   sMMMh     .odNMMMMNd+`   `+dNMMMMNdo.    \033[33m");        
  $display("                     .o---yMMdsdo------------------------:s`             \033[36m MMMMNmmmdho-     dMMMdooosMMMM+      `./sdNMMMd.    `.:ohNMMMm-   \033[33m");        
  $display("                    -yo:--/hmmds:----------------//:------o              \033[34m MMMM:...        sMMMMMMMMMMMMMN-  ``     `:MMMM+ ``      -NMMMs   \033[33m");        
  $display("                   /yssy----:::-------o+-------/h/-hy:---:+              \033[34m MMMM:          /MMMN:------hMMMd  +dy+:::/yMMMN- :my+:::/sMMMM/   \033[33m");        
  $display("                  :ysssh:------//////++/-------sMdyNMo---o.              \033[35m MMMM:         /mMMMs       .NMMMs  NMMMMMMMMmh/   NMMMMMMMMNh/    \033[33m");        
  $display("                  ossssh:-------ddddmmmds/:----:hmNNh:---o               \033[30m`::::`         .::::`        -:::: `-:/++++/-.     .:/++++/-.      \033[33m");        
  $display("                  /yssyo--------dhhyyhhdmmhy+:---://----+-                                                                                  ");        
  $display("                  `yss+---------hoo++oosydms----------::s    .......                                                                       ");        
  $display("                   :+-----------y+++++++oho--------:+sssy.://:::://+o.                                                                      ");        
  $display("                    //----------y++++++os/--------+yssssy/:--------:/s-                                                                     ");        
  $display("              ..:::::s+//:::----+s+++ooo:--------+yssssy:-----------++                                                                      ");        
  $display("            ://::------::///+/:--+soo+:----------ssssys/---------:o+s.                                                                     ");        
  $display("          .+:----------------/++/:---------------:sys+----------:o/////////::::-...                                                         ");        
  $display("          o---------------------oo::----------::/+//---------::o+--------------:/ohdhyo/-.                                                 ");        
  $display("          o---------------------/s+////:----:://:---------::/+h/------------------:oNMMMMNmhs+:.                                            ");        
  $display("          -+:::::--------------:s+-:::-----------------:://++:s--::------------::://sMMMMMMMMMMNds                                          ");        
  $display("           .+++/////////////+++s/:------------------:://+++- :+--////::------/ydmNNMMMMMMMMMMMMMMmo                                         ");        
  $display("             ./+oo+++oooo++/:---------------------:///++/-   o--:///////::----sNMMMMMMMMMMMMMMMmo                                           ");        
  $display("                o::::::--------------------------:/+++:`    .o--////////////:--+mMMMMMMMMMMMMmo                                             ");        
  $display("               :+--------------------------------/so.       +:-:////+++++///++//+mMMMMMMMMMmo                                               ");        
  $display("              .s----------------------------------+: ````` `s--////o:.-:/+syddmNMMMMMMMMMmo                                                 ");        
  $display("              o:----------------------------------s. :s+/////--//+o-        -:+shmNNMMMNs                                                   ");        
  $display("             //-----------------------------------s` .s///:---:/+o.                -/+o                                                     ");        
  $display("            .o------------------------------------o.  y///+//:/+o                                                                           ");        
  $display("            o-------------------------------------:/  o+//s//+++                                                                            ");        
  $display("           //--------------------------------------s+/o+//s                                                                                 ");        
  $display("          -+---------------------------------------:y++///s                                                                                 ");        
  $display("          o-----------------------------------------oo/+++o                                                                                 ");        
  $display("          s-----------------------------------------:s                                                                                    ");        
  $display("          o-:::::------------------:::::-------------o                                                                                      ");        
  $display("           +//////////::::::://///////////////:::----o                                                                                      ");        
  $display("           :soo+///////////+++oooooo+/////////////:-//                                                                                      ");        
  $display("       -/os/--:++/+ooo:::---..:://+ooooo++///////++so-                                                                                      ");        
  $display("      syyooo+o++//::-                   -::/yoooo+/:::+s/.                                                                                  ");        
  $display("                                             -::::///:++sys:                                                                                ");        
  $display("                                                     .:::/o+  \033[37m                                                                              ");	
  $display(" 																															");

$display ("----------------------------------------------------------------------------------------------------------------------");
$display ("                                                  Congratulations!                						            ");
$display ("----------------------------------------------------------------------------------------------------------------------");
$finish;	
end endtask


endmodule