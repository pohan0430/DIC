//==============================================
//==============================================				
//	Author	:	Wei Lu																		
//----------------------------------------------
//												
//	File Name		:	Adder_4bit.v					
//	Module Name		:	Adder_4bit					
//	Release version	:	v1.0					
//												
//----------------------------------------------								
//----------------------------------------------											
//	Input	:   A,
//				B,												
//	Output	:	Output,					
//==============================================
//==============================================
module Adder_4bit(
    //Input Port
	A,	
	B,
    //Output Port
	Output
    );

//---------------------------------------------------------------------
//   PORT DECLARATION
//---------------------------------------------------------------------
input [3:0]A;
input [3:0]B;

output wire [4:0]Output;


assign Output = A + B;


endmodule