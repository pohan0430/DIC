//==============================================
//==============================================				
//	Author	:	Wei Lu																		
//----------------------------------------------
//												
//	File Name		:	Adder_4bit.v					
//	Module Name		:	Adder_4bit					
//	Release version	:	v1.0					
//												
//----------------------------------------------								
//----------------------------------------------											
//	Input	:   A,
//				B,												
//	Output	:	Output,					
//==============================================
//==============================================
module Adder_4bit(
    //Input Port
	A,	
	B,
    //Output Port
	sum,carry
    );

//---------------------------------------------------------------------
//   PORT DECLARATION
//---------------------------------------------------------------------
input [3:0]A;
input [3:0]B;

output wire [3:0]sum;
output wire carry;


assign {carry,sum} = A + B;


endmodule
